module decoder_5to32
(
    input [4:0] IN,
    output reg [31:0] OUT
);

always @(*) begin
    case(IN)
        5'd0:  OUT = 32'b00000000000000000000000000000001;
        5'd1:  OUT = 32'b00000000000000000000000000000010;
        5'd2:  OUT = 32'b00000000000000000000000000000100;
        5'd3:  OUT = 32'b00000000000000000000000000001000;
        5'd4:  OUT = 32'b00000000000000000000000000010000;
        5'd5:  OUT = 32'b00000000000000000000000000100000;
        5'd6:  OUT = 32'b00000000000000000000000001000000;
        5'd7:  OUT = 32'b00000000000000000000000010000000;
        5'd8:  OUT = 32'b00000000000000000000000100000000;
        5'd9:  OUT = 32'b00000000000000000000001000000000;
        5'd10: OUT = 32'b00000000000000000000010000000000;
        5'd11: OUT = 32'b00000000000000000000100000000000;
        5'd12: OUT = 32'b00000000000000000001000000000000;
        5'd13: OUT = 32'b00000000000000000010000000000000;
        5'd14: OUT = 32'b00000000000000000100000000000000;
        5'd15: OUT = 32'b00000000000000001000000000000000;
        5'd16: OUT = 32'b00000000000000010000000000000000;
        5'd17: OUT = 32'b00000000000000100000000000000000;
        5'd18: OUT = 32'b00000000000001000000000000000000;
        5'd19: OUT = 32'b00000000000010000000000000000000;
        5'd20: OUT = 32'b00000000000100000000000000000000;
        5'd21: OUT = 32'b00000000001000000000000000000000;
        5'd22: OUT = 32'b00000000010000000000000000000000;
        5'd23: OUT = 32'b00000000100000000000000000000000;
        5'd24: OUT = 32'b00000001000000000000000000000000;
        5'd25: OUT = 32'b00000010000000000000000000000000;
        5'd26: OUT = 32'b00000100000000000000000000000000;
        5'd27: OUT = 32'b00001000000000000000000000000000;
        5'd28: OUT = 32'b00010000000000000000000000000000;
        5'd29: OUT = 32'b00100000000000000000000000000000;
        5'd30: OUT = 32'b01000000000000000000000000000000;
        5'd31: OUT = 32'b10000000000000000000000000000000;
        default: OUT = 32'b0;
    endcase
end

endmodule
